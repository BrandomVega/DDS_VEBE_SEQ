LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DETECTOR IS 
	PORT( CLK :IN STD_LOGIC;
	CLR: IN STD_LOGIC;						
	ENB: IN STD_LOGIC;
	ENTRADA: IN STD_LOGIC_VECTOR(6 DOWNTO 0);
	SALIDA: OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END DETECTOR;

ARCHITECTURE COMPORTAMENTAL OF DETECTOR IS 
TYPE ESTADOS IS(A, B, C, D, E, F, G);		  
attribute ENUM_ENCODING: STRING;
ATTRIBUTE enum_encoding OF ESTADOS: TYPE IS
"0000" & --A--	  
"0001" & --B--
"0011" & --C--
"0010" & --D--
"0110" & --E--
"0111" & --F--
"1111" ; --G--
SIGNAL EDO, NEXT_EDO: ESTADOS;
SIGNAL AUX_ENTRADA: STD_LOGIC_VECTOR(6 DOWNTO 0);
SIGNAL AUX_SALIDA: STD_LOGIC;
BEGIN

PROCESS (CLR, CLK, ENB)
BEGIN 
	IF(CLR = '1') THEN
		EDO <= A;						   
	ELSIF(ENB = '1') THEN
	   EDO <= EDO;						   
	ELSIF(CLK'EVENT AND CLK = '1') THEN
		EDO <= NEXT_EDO;
	END IF;
END PROCESS;	   

PROCESS(CLK, CLR) BEGIN
		IF (CLR ='1') THEN
			AUX_ENTRADA <= (OTHERS => '0');
		ELSIF (ENB = '1') THEN 
			AUX_ENTRADA <= ENTRADA;
		ELSIF (CLK'EVENT AND CLK = '1') THEN 
			AUX_ENTRADA(5 DOWNTO 0) <= AUX_ENTRADA(6 DOWNTO 1);
			AUX_ENTRADA(6) <= '0';
		END IF;
END PROCESS;
AUX_SALIDA <= AUX_ENTRADA(0);

PROCESS (AUX_SALIDA, EDO)
BEGIN 
	CASE EDO IS WHEN 
		A => IF AUX_SALIDA = '0' THEN
			NEXT_EDO <= C;
		ELSIF AUX_SALIDA = '1' THEN
			NEXT_EDO <= B;
		END IF;
		WHEN
		B => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF AUX_SALIDA = '1' THEN
			NEXT_EDO  <= F;
		END IF;	
		WHEN
		C => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= D;
		ELSIF AUX_SALIDA ='1' THEN
			NEXT_EDO <= B;
		END IF;
		WHEN
		D => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= E;
		ELSIF AUX_SALIDA ='1' THEN
			NEXT_EDO <= B;
		END IF;			 
		WHEN
		E => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= E;
		ELSIF AUX_SALIDA ='1' THEN
			NEXT_EDO <= B;
		END IF;			  
		WHEN
		F => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF AUX_SALIDA ='1' THEN
			NEXT_EDO <= G;
		END IF;			  
		WHEN
		G => IF AUX_SALIDA = '0' THEN 
			NEXT_EDO <= C;
		ELSIF AUX_SALIDA ='1' THEN
			NEXT_EDO <= G;
		END IF;		   
		WHEN OTHERS => NULL;
	END CASE;
END PROCESS;
--A B C D E F G--
SALIDA <= "0110000" WHEN (EDO = C AND AUX_SALIDA = '0') ELSE--A--
	"0110000" WHEN (EDO = B AND AUX_SALIDA = '1' ) ELSE 
	"0110000" WHEN (EDO = C AND AUX_SALIDA = '0') ELSE --B--
	"0110000" WHEN (EDO = F AND AUX_SALIDA = '1' ) ELSE
	"0110000" WHEN (EDO = D AND AUX_SALIDA = '0') ELSE --C--
	"0110000" WHEN (EDO = B AND AUX_SALIDA = '1' ) ELSE
	"0001001" WHEN (EDO = E AND AUX_SALIDA = '0') ELSE	--D--
	"0110000" WHEN (EDO = B AND AUX_SALIDA = '1' ) ELSE 
	"0001001" WHEN (EDO = E AND AUX_SALIDA = '0') ELSE	 --E-
	"0110000" WHEN (EDO = B AND AUX_SALIDA = '1' ) ELSE
	"0110000" WHEN (EDO = C AND AUX_SALIDA = '0') ELSE	--F--
	"0001001" WHEN (EDO = G AND AUX_SALIDA = '1' ) ELSE
	"0110000" WHEN (EDO = B AND AUX_SALIDA = '0') ELSE	--G
	"0001001" WHEN (EDO = G AND AUX_SALIDA = '1' ) ELSE   
	"0110000";
END COMPORTAMENTAL;
		
	

		
		

