

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;


ENTITY SIPO IS
	PORT(
	CLK, CLR: IN STD_LOGIC;
	Q: INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);	   
	D: IN STD_LOGIC);
END ENTITY;

ARCHITECTURE SIPO OF SIPO IS

BEGIN
	PROCESS(CLK, CLR) BEGIN		  
		IF(CLR = '1')THEN
			Q <= (OTHERS => '0');
		ELSIF(CLK'EVENT AND CLK='1')THEN
		  	Q(3) <= D; 
			Q(2 DOWNTO 0) <= Q(3 DOWNTO 1);
		END IF;
	END PROCESS;
END ARCHITECTURE;