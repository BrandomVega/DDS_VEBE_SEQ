

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY SISO IS
	PORT(	   
		CLK, CLR, D: IN STD_LOGIC;
		Q4: OUT STD_LOGIC	
	);
END ENTITY;
	
ARCHITECTURE SISO OF SISO IS
SIGNAL QAUX: STD_LOGIC_VECTOR(3 DOWNTO 1);
BEGIN			
	PROCESS(CLR, CLK) BEGIN		
		IF(CLR='1')THEN
			Q4<='0';
			QAUX<=(OTHERS=>'0'); 
		ELSIF(CLK'EVENT AND CLK='1')THEN
			QAUX(1)<=D;
			QAUX(3 DOWNTO 2) <= QAUX(2 DOWNTO 1);
			Q4 <= QAUX(3);
		END IF;
	END PROCESS;
END ARCHITECTURE;