LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;		   

ENTITY PISO IS
	PORT(	   
		CLK, CLR, SHIFTLOAD: IN STD_LOGIC;
		D: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		QN: OUT STD_LOGIC	
	);
END ENTITY;
	
ARCHITECTURE PISO OF PISO IS
SIGNAL QAUX: STD_LOGIC_VECTOR(3 DOWNTO 0);
BEGIN			
	PROCESS(CLR, CLK) BEGIN		
		IF(CLR='1')THEN
			QAUX <= (OTHERS => '0');
		ELSIF(CLK'EVENT AND CLK='1')THEN 
			IF(SHIFTLOAD = '1')THEN
				QAUX<=D;	
			ELSE
				QAUX(2 DOWNTO 0) <= QAUX(3 DOWNTO 1);  
				QAUX(3)<='0';
			END IF;	   
		END IF;	
	END PROCESS;   
	QN <= QAUX(0);
END ARCHITECTURE;


